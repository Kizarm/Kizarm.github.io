.title lambda oscilator
.global gnd
c1 out 0 1.5u ic=5
r1 out net-_r1-pad2_ 100m
xr1 net-_v1-pad1_ drv lambda
xl1 0 net-_r1-pad2_ drv p1s3
v1 net-_v1-pad1_ 0 2.5
.model pmbfj177 pjf vto=-1.8000e+000 beta=3.37432e-003 lambda=2.41676e-002 rd=1.45880e+000 rs=1.45880e+000 is=7.27555e-016 cgs=8.90000e-012 cgd=1.02500e-011 pb=6.94243e-001 fc=5.00000e-001
.model pmbfj112 njf vto=-2.3303e+000 beta=5.97264e-003 lambda=2.31986e-002 rd=2.29075e+000 rs=2.29075e+000 is=8.87988e-016 cgs=1.05000e-011 cgd=1.20000e-011 pb=6.09944e-001 fc=5.00000e-001
.subckt p1s3 1 2 3
l01 3 2 10m
l02 1 3 1m
k01 l01 l02 1
.ends p1s3
.subckt lambda a b
j01 a b c pmbfj112
j02 c a b pmbfj177
.ends lambda
vxx1 out /out 0
vxx2 drv /drv 0
.tran 1u 10m uic
.end
