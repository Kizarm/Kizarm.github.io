.title delic
.global gnd
.model qbc847 npn is=1.822e-14 nf=0.9932 ise=2.894e-16 ne=1.4 bf=324.4 ikf=0.109 vaf=82 nr=0.9931 isc=9.982e-12 nc=1.763 br=8.29 ikr=0.09 var=17.9 rb=10 irb=5e-06 rbm=5 re=0.649 rc=0.7014 xtb=0 eg=1.11 xti=3 cje=1.244e-11 vje=0.7579 mje=0.3656 tf=4.908e-10 xtf=9.51 vtf=2.927 itf=0.3131 ptf=0 cjc=3.347e-12 vjc=0.5463 mjc=0.391 xcjc=0.6193 tr=9e-08 cjs=0 vjs=0.75 mjs=0.333 fc=0.979
v2 in 0 pulse(1.2 2.8 0 1u 1u 4u 10u ) dc=0
r1 in net-_q1-pad1_ 8k
q2 t2 net-_q1-pad1_ net-_q2-pad3_ qbc847
q1 net-_q1-pad1_ t2 net-_q1-pad3_ qbc847
r2 in t2 8k
r3 net-_r10-pad1_ net-_q3-pad1_ 1k
q4 t1 net-_q1-pad3_ 0 qbc847
q3 net-_q3-pad1_ net-_q2-pad3_ 0 qbc847
r4 net-_r10-pad1_ t1 1k
r5 net-_q1-pad3_ net-_q3-pad1_ 4k
r6 t1 net-_q2-pad3_ 4k
v1 net-_r10-pad1_ 0 6
r8 t1 net-_q5-pad1_ 8k
q6 t4 net-_q5-pad1_ net-_q6-pad3_ qbc847
q5 net-_q5-pad1_ t4 net-_q5-pad3_ qbc847
r9 t1 t4 8k
r7 net-_r10-pad1_ net-_q7-pad1_ 1k
q8 t3 net-_q5-pad3_ 0 qbc847
q7 net-_q7-pad1_ net-_q6-pad3_ 0 qbc847
r10 net-_r10-pad1_ t3 1k
r11 net-_q5-pad3_ net-_q7-pad1_ 4k
r12 t3 net-_q6-pad3_ 4k
**************************
vx0 in /in 0
vx1 t1 /t1 0
vx2 t2 /t2 0
vx3 t3 /t3 0
vx4 t4 /t4 0
.tran 10n 100u
.end
