.title bistable cmos
.subckt SXN 1 2 3
M01 1 2 3 3 MMN
C01 2 3 100p
.MODEL MMN NMOS LEVEL=1 VTO=1 KP=8m
.ends SXN
.subckt SXP 1 2 3
M02 1 2 3 3 MMP
C02 2 3 100p
.MODEL MMP PMOS LEVEL=1 VTO=-1.1 KP=8m
.ends SXP
*********************
V1  VCC 0 5		
XQ1 /OUT /MID VCC SXP
XQ2 /OUT /MID 0   SXN
XQ3 /MID /INP VCC SXP
XQ4 /MID /INP 0   SXN
C1  /INP /OUT 5n IC=2
R1  /MID /INP 10k
*********************
.tran 100n 500u uic
.end
